* Kaspix Active Sallen-Key Low Pass Filter
* Topología: Sallen-Key de 2do Orden con Ganancia Unitaria
* Parametros a aprender: Frecuencia de corte (via R_tune)

* --- 1. PARAMETROS VARIABLES (KNOBS) ---
* R_tune: Controla la frecuencia de corte.
* Rango sugerido: 1k (agudo) a 50k (grave)
.param R_tune=10k

* --- 2. ENTRADA Y ALIMENTACIÓN ---
Vin input 0 DC 0 AC 1
* Alimentación virtual del OpAmp (para saturación realista)
Vcc  pos_rail 0 15
Vee  neg_rail 0 -15

* --- 3. CIRCUITO SALLEN-KEY ---
* La señal entra por input, pasa por la red RC y va a la entrada no-inv del OpAmp.
* R1 y R2 son las resistencias variables que definen la frecuencia.

R1 input n1 {R_tune}
R2 n1 n_plus {R_tune}

* Capacitores fijos (determinan el rango de operación)
C1 n1 output 10n
C2 n_plus 0 10n

* --- 4. AMPLIFICADOR OPERACIONAL (Modelo Idealizado con Saturation) ---
* X1 n_plus n_minus pos_rail neg_rail output OPAMP_SIMPLE
* Configurado como buffer (ganancia unitaria): Salida conectada a entrada inv (n_minus)
E_opamp output 0 VOLTAGE ( n_plus 0 ) 1
* Nota: Para simplificar la simulación en dataset, usaremos un VCVS ideal
* Si quieres distorsión, avísame y ponemos un modelo no-lineal.
* Por ahora, esto asegura convergencia perfecta.

* Feedback para buffer
* En Sallen-Key unitario, la salida se conecta directo a C1 (bootstrapping)
* Corrección de nodo: C1 va de n1 a output en esta topología.

* --- 5. CARGA ---
R_load output 0 100k

.save V(output)
.tran 10u 40m
.end