* Kaspix Standardized High-Pass Filter (HPF)
* Propósito: Filtro de primer orden para eliminación de graves.

.param R_gain=10k    ; Resistencia a tierra (1k - 100k)
.param C_hp=100n     ; Capacitor en serie (10n - 1u)

* Entrada y Fuente
Vin input 0 DC 0 AC 1

* Circuito CR
C1 input output {C_hp}
R1 output 0 {R_gain}

* Carga
RLoad output 0 1Meg

.save V(output)
.end